

 
 
 

 



window new WaveWindow  -name  "Waves for BMG Example Design"
waveform  using  "Waves for BMG Example Design"

      waveform add -signals /Win_RAM_tb/status
      waveform add -signals /Win_RAM_tb/Win_RAM_synth_inst/bmg_port/CLKA
      waveform add -signals /Win_RAM_tb/Win_RAM_synth_inst/bmg_port/ADDRA
      waveform add -signals /Win_RAM_tb/Win_RAM_synth_inst/bmg_port/DINA
      waveform add -signals /Win_RAM_tb/Win_RAM_synth_inst/bmg_port/WEA
      waveform add -signals /Win_RAM_tb/Win_RAM_synth_inst/bmg_port/DOUTA

console submit -using simulator -wait no "run"
